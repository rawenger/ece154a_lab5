// lab 5 controller FSM testbench
module controller_tb();

endmodule